module AudPlayer(
    input i_rst_n,
    input i_bclk,
    input i_daclrck,
    input i_en,
    input i_dac_data,
    output o_aud_dacdat
);

endmodule